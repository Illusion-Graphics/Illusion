`ifndef __DEFINES_SVH
`define __DEFINES_SVH

typedef enum [15:0] {
	COMMAND_OP_FLOAT_INT = 16'h0001,
	COMMAND_OP_INT_FLOAT = 16'h0002
} Commands;

`endif // __DEFINES_SVH
